/////////////////////////////////////////////////////
//
//  // HEADER //
//
//  FILE NAME = axi_s_defines.svh
//  ENGINEER  = Muskan
//  VERSION   = 1.0 
//  DESCRIPTION = contains all macro 
//
/////////////////////////////////////////////////////

`ifndef AXI_S_DEFINES
`define AXI_S_DEFINES

 `define DATA_WIDTH;
 `define ADD_WIDTH;

`endif
