/////////////////////////////////////////////////////
//
//  // HEADER //
//
//  FILE NAME = axi_m_defines.svh
//  ENGINEER  = Muskan
//  VERSION   = 1.0 
//  DESCRIPTION = contains all macro 
//
/////////////////////////////////////////////////////

`ifndef AXI_M_DEFINES
`define AXI_M_DEFINES

 `define DATA_WIDTH;
 `define ADD_WIDTH;

`endif
